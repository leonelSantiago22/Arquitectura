

library IEEE;
use IEEE.STD_LOGIC_1164.all;



entity burbuja_instruccion is
	 port(
		 salida : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end burbuja_instruccion;

--}} End of automatically maintained section

architecture burbuja_instruccion of burbuja_instruccion is
begin
	
		salida<= x"00000000";
	 -- enter your statements here --

end burbuja_instruccion;
